------------------------------------------------------
-- LogiBLOX ROM Module "rom64x16"
-- Created by LogiBLOX version C.16
--    on Fri May 27 02:20:32 2011
-- Attributes 
--    MODTYPE = ROM
--    BUS_WIDTH = 16
--    DEPTH = 128
--    MEMFILE = rom
--    TRIM = FALSE
--    STYLE = MAX_SPEED
--    USE_RPM = FALSE
------------------------------------------------------
-- This is a behaviorial model only and cannot be synthesized.
------------------------------------------------------
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
LIBRARY logiblox;
USE logiblox.mvlutil.ALL;
USE logiblox.mvlarith.ALL;
USE logiblox.logiblox.ALL;

ENTITY rom64x16 IS
  PORT(
    A: IN std_logic_vector(6 DOWNTO 0);
    DO: OUT std_logic_vector(15 DOWNTO 0));
END rom64x16;

ARCHITECTURE sim OF rom64x16 IS
  SIGNAL START_PULSE: std_logic := '1';
  TYPE mem_data IS ARRAY (127 DOWNTO 0) OF std_logic_vector(15 DOWNTO 0);
BEGIN
  PROCESS
  VARIABLE VD: mem_data;
  VARIABLE first_time: BOOLEAN := TRUE;
  BEGIN
    IF (first_time) THEN
      VD(0) := ('0','1','0','0','1','0','0','1','0','0','1','0','0','0','0','0');
      VD(1) := ('0','1','0','0','1','0','1','0','0','1','0','0','0','0','0','0');
      VD(2) := ('0','1','0','0','1','0','1','1','0','1','1','0','0','0','0','0');
      VD(3) := ('0','1','0','0','1','1','0','0','1','0','0','0','0','0','0','0');
      VD(4) := ('0','1','0','0','1','1','0','1','1','0','1','0','0','0','0','0');
      VD(5) := ('0','1','0','0','1','1','1','0','1','1','0','0','0','0','0','0');
      VD(6) := ('0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0');
      VD(7) := ('0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','1');
      VD(8) := ('1','1','0','0','1','1','1','1','0','1','0','1','0','1','1','0');
      VD(9) := ('0','1','0','0','1','1','1','1','1','1','1','0','0','0','0','0');
      VD(10) := ('0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0');
      VD(11) := ('1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','1');
      VD(12) := ('1','1','0','0','1','1','1','1','0','1','0','1','0','1','1','1');
      VD(13) := ('0','1','0','0','1','1','1','1','1','1','1','0','0','0','0','0');
      VD(14) := ('0','0','0','0','0','0','0','0','0','1','1','1','0','0','0','0');
      VD(15) := ('1','1','1','1','1','1','1','1','1','1','1','1','1','0','1','0');
      VD(16) := ('1','1','0','0','1','1','1','1','0','1','0','1','1','0','0','0');
      VD(17) := ('0','1','0','0','1','1','1','1','1','1','1','0','0','0','0','0');
      VD(18) := ('0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0');
      VD(19) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1');
      VD(20) := ('1','1','0','0','1','1','1','1','0','1','0','1','1','0','0','1');
      VD(21) := ('0','1','0','0','1','1','1','1','1','1','1','0','0','0','0','0');
      VD(22) := ('0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0');
      VD(23) := ('0','0','0','0','0','0','0','0','0','0','0','1','0','1','1','1');
      VD(24) := ('1','1','0','0','1','1','1','1','0','1','0','1','1','0','1','0');
      VD(25) := ('0','1','0','0','1','1','1','1','1','1','1','0','0','0','0','0');
      VD(26) := ('0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0');
      VD(27) := ('1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1');
      VD(28) := ('1','1','0','0','1','1','1','1','0','1','0','1','1','0','1','1');
      VD(29) := ('0','1','0','0','1','1','1','1','1','1','1','0','0','0','0','0');
      VD(30) := ('0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0');
      VD(31) := ('1','1','1','1','1','1','1','1','1','1','1','1','1','1','0','0');
      VD(32) := ('1','1','0','0','1','1','1','1','0','1','0','1','1','1','0','0');
      VD(33) := ('0','1','0','0','1','1','1','1','1','1','1','0','0','0','0','0');
      VD(34) := ('0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0');
      VD(35) := ('1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1');
      VD(36) := ('1','1','0','0','1','1','1','1','0','1','0','1','1','1','0','1');
      VD(37) := ('0','1','0','0','1','1','1','1','1','1','1','0','0','0','0','0');
      VD(38) := ('0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0');
      VD(39) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','1','0','0');
      VD(40) := ('1','1','0','0','1','1','1','1','0','1','0','1','1','1','1','0');
      VD(41) := ('0','1','0','0','1','1','1','1','1','1','1','0','0','0','0','0');
      VD(42) := ('0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0');
      VD(43) := ('0','0','0','0','0','0','0','0','0','0','1','1','0','1','1','0');
      VD(44) := ('1','1','0','0','1','1','1','1','0','1','0','1','1','1','1','1');
      VD(45) := ('0','1','0','0','1','1','1','1','1','1','1','0','0','0','0','0');
      VD(46) := ('0','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0');
      VD(47) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1');
      VD(48) := ('1','1','0','0','0','0','1','0','0','0','1','1','1','1','1','0');
      VD(49) := ('1','1','0','0','0','0','1','1','0','0','1','1','1','1','1','1');
      VD(50) := ('0','0','0','0','1','0','1','1','0','0','0','0','0','0','0','0');
      VD(51) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1');
      VD(52) := ('1','1','0','0','0','1','0','0','0','0','1','1','1','1','1','1');
      VD(53) := ('1','1','0','0','0','1','0','0','0','0','1','1','1','1','1','0');
      VD(54) := ('1','0','0','0','0','1','0','1','0','0','1','1','1','1','1','1');
      VD(55) := ('0','1','0','0','0','1','0','0','0','1','0','0','0','0','0','0');
      VD(56) := ('1','1','0','0','1','1','0','0','0','0','1','1','1','1','1','1');
      VD(57) := ('1','0','0','0','1','1','0','1','0','0','1','1','1','1','1','1');
      VD(58) := ('1','1','1','0','1','1','1','1','1','0','1','0','0','0','0','0');
      VD(59) := ('0','0','0','0','0','0','0','0','0','0','1','1','1','1','1','0');
      VD(60) := ('0','1','0','0','0','0','0','1','1','0','1','0','0','0','0','0');
      VD(61) := ('1','1','1','0','0','0','0','0','0','1','0','0','0','0','0','0');
      VD(62) := ('0','1','0','0','1','0','0','1','1','0','1','0','0','0','0','0');
      VD(63) := ('1','1','1','0','0','0','0','0','0','1','0','0','0','0','0','0');
      VD(64) := ('0','1','0','0','1','1','0','0','0','1','1','0','0','0','0','0');
      VD(65) := ('1','1','0','0','1','1','0','0','0','0','1','1','1','1','1','1');
      VD(66) := ('0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0');
      VD(67) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1');
      VD(68) := ('1','1','1','0','1','1','1','1','1','1','0','0','0','0','0','0');
      VD(69) := ('0','0','0','0','0','0','0','0','0','1','0','0','0','1','1','1');
      VD(70) := ('1','1','1','0','0','0','0','0','0','0','1','1','0','1','1','0');
      VD(71) := ('1','1','0','0','1','0','0','1','0','1','0','0','0','0','0','0');
      VD(72) := ('1','1','0','1','1','0','0','1','0','0','0','0','0','0','0','0');
      VD(73) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(74) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(75) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(76) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(77) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(78) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(79) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(80) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(81) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(82) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(83) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(84) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(85) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(86) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(87) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(88) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(89) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(90) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(91) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(92) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(93) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(94) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(95) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(96) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(97) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(98) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(99) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(100) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(101) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(102) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(103) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(104) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(105) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(106) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(107) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(108) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(109) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(110) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(111) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(112) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(113) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(114) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(115) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(116) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(117) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(118) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(119) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(120) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(121) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(122) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(123) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(124) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(125) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(126) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(127) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      first_time := FALSE;
    END IF;
    IF (mvlvec_not01(A)) THEN
      DO <= ('X','X','X','X','X','X','X','X','X','X','X','X','X','X','X','X');
    ELSE
      DO <= VD(mvlvec2int(A));
    END IF;
      WAIT ON A, START_PULSE;
  END PROCESS;
END sim;
