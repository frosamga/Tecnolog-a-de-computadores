------------------------------------------------------
-- LogiBLOX SYNC_RAM Module "ram256x16"
-- Created by LogiBLOX version C.16
--    on Thu Feb 18 13:10:44 2010
-- Attributes 
--    MODTYPE = SYNC_RAM
--    BUS_WIDTH = 16
--    DEPTH = 256
--    STYLE = MAX_SPEED
--    USE_RPM = FALSE
------------------------------------------------------
-- This is a behaviorial model only and cannot be synthesized.
------------------------------------------------------
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
LIBRARY logiblox;
USE logiblox.mvlutil.ALL;
USE logiblox.mvlarith.ALL;
USE logiblox.logiblox.ALL;

ENTITY ram256x16 IS
  PORT(
    A: IN std_logic_vector(7 DOWNTO 0);
    DO: OUT std_logic_vector(15 DOWNTO 0);
    DI: IN std_logic_vector(15 DOWNTO 0);
    WR_EN: IN std_logic;
    WR_CLK: IN std_logic);
END ram256x16;

ARCHITECTURE sim OF ram256x16 IS
  SIGNAL START_PULSE: std_logic := '1';
  TYPE mem_data IS ARRAY (255 DOWNTO 0) OF std_logic_vector(15 DOWNTO 0);
BEGIN
  PROCESS
  VARIABLE VD: mem_data;
  VARIABLE first_time: BOOLEAN := TRUE;
  BEGIN
    IF (first_time) THEN
      VD(0) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(1) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(2) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(3) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(4) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(5) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(6) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(7) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(8) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(9) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(10) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(11) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(12) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(13) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(14) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(15) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(16) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(17) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(18) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(19) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(20) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(21) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(22) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(23) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(24) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(25) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(26) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(27) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(28) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(29) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(30) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(31) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(32) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(33) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(34) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(35) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(36) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(37) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(38) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(39) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(40) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(41) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(42) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(43) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(44) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(45) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(46) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(47) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(48) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(49) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(50) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(51) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(52) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(53) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(54) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(55) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(56) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(57) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(58) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(59) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(60) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(61) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(62) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(63) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(64) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(65) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(66) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(67) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(68) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(69) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(70) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(71) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(72) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(73) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(74) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(75) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(76) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(77) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(78) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(79) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(80) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(81) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(82) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(83) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(84) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(85) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(86) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(87) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(88) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(89) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(90) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(91) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(92) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(93) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(94) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(95) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(96) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(97) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(98) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(99) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(100) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(101) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(102) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(103) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(104) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(105) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(106) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(107) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(108) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(109) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(110) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(111) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(112) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(113) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(114) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(115) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(116) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(117) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(118) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(119) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(120) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(121) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(122) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(123) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(124) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(125) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(126) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(127) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(128) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(129) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(130) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(131) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(132) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(133) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(134) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(135) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(136) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(137) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(138) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(139) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(140) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(141) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(142) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(143) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(144) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(145) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(146) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(147) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(148) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(149) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(150) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(151) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(152) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(153) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(154) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(155) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(156) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(157) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(158) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(159) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(160) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(161) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(162) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(163) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(164) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(165) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(166) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(167) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(168) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(169) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(170) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(171) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(172) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(173) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(174) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(175) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(176) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(177) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(178) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(179) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(180) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(181) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(182) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(183) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(184) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(185) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(186) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(187) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(188) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(189) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(190) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(191) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(192) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(193) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(194) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(195) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(196) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(197) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(198) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(199) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(200) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(201) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(202) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(203) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(204) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(205) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(206) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(207) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(208) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(209) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(210) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(211) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(212) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(213) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(214) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(215) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(216) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(217) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(218) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(219) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(220) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(221) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(222) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(223) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(224) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(225) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(226) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(227) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(228) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(229) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(230) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(231) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(232) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(233) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(234) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(235) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(236) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(237) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(238) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(239) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(240) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(241) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(242) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(243) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(244) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(245) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(246) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(247) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(248) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(249) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(250) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(251) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(252) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(253) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(254) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      VD(255) := ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
      first_time := FALSE;
    END IF;
    IF (WR_CLK'EVENT AND stdbit2mvl(WR_CLK)='1' AND stdbit2mvl(WR_CLK'LAST_VALUE)='0')
    AND (WR_EN='1') AND (NOT mvlvec_not01(A)) THEN
      VD(mvlvec2int(A)) := stdvec2mvl(DI);
    END IF;
    IF (mvlvec_not01(A) OR
       (stdbit2mvl(WR_CLK) = 'X')
       OR (WR_CLK'EVENT AND stdbit2mvl(WR_CLK)='1' AND stdbit2mvl(WR_CLK'LAST_VALUE)='0'
           AND stdbit2mvl(WR_EN) = 'X' )
      ) THEN
        DO <= ('X','X','X','X','X','X','X','X','X','X','X','X','X','X','X','X');
    ELSE
      DO <= VD(mvlvec2int(A));
    END IF;
      WAIT ON A, DI, WR_EN, WR_CLK, START_PULSE;
  END PROCESS;
END sim;
